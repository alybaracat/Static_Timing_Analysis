`timescale 1ns/1ns

module simple_design1(a,b,y);
input a,b;
output y;

assign y = a & b;

endmodule
